module led_blinking(led);
	output[7:0] led;
			assign led=8'b10101010;
endmodule